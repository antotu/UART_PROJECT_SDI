library ieee;
use ieee.std_logic_1164.all;


entity CU_RX is 
port (
CLK : IN STD_LOGIC;

-- INPUT
EN_RX : IN STD_LOGIC;
ERROR_STATUS : IN STD_LOGIC;
START : IN STD_LOGIC;
TC_TIME_SAMPLE : IN STD_LOGIC;
TC_8_SAMPLES : IN STD_LOGIC;
TC_4_SAMPLES : IN STD_LOGIC;
TC_READ_ALL : IN STD_LOGIC;
TC_TIME_NOP : IN STD_LOGIC;

-- OUTPUT
CLEAR_DOUT : OUT STD_LOGIC;
LD_SHIFT_R8 : OUT STD_LOGIC;
CLEAR_R8 : OUT STD_LOGIC;
MUX_SEL_STOP_BIT : OUT STD_LOGIC;
LD_ERROR : OUT STD_LOGIC;
CLEAR_ERROR : OUT STD_LOGIC;
CLEAR_BUSY : OUT STD_LOGIC;
LD_BUSY : OUT STD_LOGIC;
LD_SHIFT_DOUT : OUT STD_LOGIC;
EN_CNT_TIME_SAMPLES : OUT STD_LOGIC;
CLEAR_CNT_TIME_SAMPLES : OUT STD_LOGIC;
EN_CNT_8_SAMPLES : OUT STD_LOGIC;
CLEAR_CNT_8_SAMPLES : OUT STD_LOGIC;
EN_CNT_SYMBOL : OUT STD_LOGIC;
CLEAR_CNT_SYMBOL : OUT STD_LOGIC;
CLEAR_DONE : OUT STD_LOGIC;
LD_DONE : OUT STD_LOGIC;

EN_CNT_TIME_NOP : OUT STD_LOGIC;
CLEAR_CNT_TIME_NOP : OUT STD_LOGIC

);
 end CU_RX;

architecture beh of CU_RX is

type STATE_TYPE is (RESET_STATE, IDLE_1, IDLE_2, STATE_AFTER_START_1, STATE_AFTER_START_2, ANALISI_SAMPLES_START_1, ANALISI_SAMPLES_START_2, LOAD_ERROR_START,
MANAGE_ERROR_START_BIT, NOP_START_SYMB, NOP_START_SYMB_END, SYMBOL_SAMPLE, SYMBOL_WAIT, EVALUATION_SYMBOLS, NOP_SYMBOL, NOP_SYMBOL_END, 
STOP_BIT_SAMPLES, STOP_BIT_WAIT,  EVALUATE_ERROR_STOP, ERROR_STOP_BIT);

SIGNAL NEXT_STATE : STATE_TYPE;
SIGNAL CURRENT_STATE : STATE_TYPE;


begin

NEXT_STATE_PROCESS: process(CURRENT_STATE, START, TC_TIME_SAMPLE, TC_8_SAMPLES, TC_4_SAMPLES, TC_READ_ALL, TC_TIME_NOP, ERROR_STATUS, EN_RX)
begin
case CURRENT_STATE is
	 WHEN RESET_STATE => if EN_RX = '1' then
				NEXT_STATE <= IDLE_1;
			else
				NEXT_STATE <= RESET_STATE;
			end if;

	WHEN IDLE_1 => NEXT_STATE <= IDLE_2;
	
	WHEN IDLE_2 => if START = '1' then
			NEXT_STATE <= STATE_AFTER_START_1;
		else
			if TC_TIME_SAMPLE = '1' then
				NEXT_STATE <= IDLE_1;
			else
				NEXT_STATE <= IDLE_2;
			end if;
		end if;
	WHEN STATE_AFTER_START_1 => NEXT_STATE <= STATE_AFTER_START_2;

	WHEN STATE_AFTER_START_2 => if TC_TIME_SAMPLE = '1' then
				NEXT_STATE <= ANALISI_SAMPLES_START_1;
				else
				NEXT_STATE <= STATE_AFTER_START_2;
				end if;
	
	WHEN ANALISI_SAMPLES_START_1 => NEXT_STATE <= ANALISI_SAMPLES_START_2;
	
	WHEN ANALISI_SAMPLES_START_2 => if TC_TIME_SAMPLE = '0' then 
					NEXT_STATE <= ANALISI_SAMPLES_START_2;
				   else
					if TC_4_SAMPLES = '0' then
					NEXT_STATE <= ANALISI_SAMPLES_START_1;
					else
					NEXT_STATE <= LOAD_ERROR_START;
					end if;
				end if;
	
	WHEN LOAD_ERROR_START => if ERROR_STATUS = '1' then
				NEXT_STATE <= MANAGE_ERROR_START_BIT;
			else
				NEXT_STATE <= NOP_START_SYMB;
			end if;
	
	
	WHEN MANAGE_ERROR_START_BIT => NEXT_STATE <= IDLE_1;

	WHEN NOP_START_SYMB => 
							if TC_TIME_NOP = '1' then
								NEXT_STATE <= NOP_START_SYMB_END;
							else
								NEXT_STATE <= NOP_START_SYMB;
							end if;
	
	WHEN NOP_START_SYMB_END => NEXT_STATE <= SYMBOL_SAMPLE;


	WHEN SYMBOL_SAMPLE => NEXT_STATE <= SYMBOL_WAIT;
	
	WHEN SYMBOL_WAIT => if TC_TIME_SAMPLE = '0' then
					NEXT_STATE <= SYMBOL_WAIT;
				
				else
					if TC_8_SAMPLES = '0' then
					NEXT_STATE <= SYMBOL_SAMPLE;
				 	else
					NEXT_STATE <= EVALUATION_SYMBOLS;
					end if;
				end if;

	WHEN EVALUATION_SYMBOLS => NEXT_STATE <= NOP_SYMBOL;

	WHEN NOP_SYMBOL => 
						if TC_TIME_NOP = '1' then
							NEXT_STATE <= NOP_SYMBOL_END;
						else
							NEXT_STATE <= NOP_SYMBOL;
						end if;

	when NOP_SYMBOL_END => 
							if TC_READ_ALL = '0' then
								NEXT_STATE <= SYMBOL_SAMPLE;
							else
								NEXT_STATE <= STOP_BIT_SAMPLES;
							end if;
	
	WHEN STOP_BIT_SAMPLES => NEXT_STATE <= STOP_BIT_WAIT;

	WHEN STOP_BIT_WAIT => if TC_8_SAMPLES = '1' then
						NEXT_STATE <= 	EVALUATE_ERROR_STOP;
					else
						if TC_TIME_SAMPLE = '0' then
							NEXT_STATE <= STOP_BIT_WAIT;
						else
						NEXT_STATE <= STOP_BIT_SAMPLES;
						end if;
					end if;
	
	WHEN EVALUATE_ERROR_STOP => if ERROR_STATUS = '1' then
				NEXT_STATE <= ERROR_STOP_BIT;
				else
				NEXT_STATE <= IDLE_2;
				end if;


	
	WHEN ERROR_STOP_BIT => NEXT_STATE <= IDLE_2;


	when others => NEXT_STATE <= RESET_STATE;


end case;

end process;


CURRENT_STATE_PROCESS : process(CLK)
begin
if CLK'EVENT AND CLK = '1' then
	if EN_RX = '0' then
		CURRENT_STATE <= RESET_STATE;
	else
		CURRENT_STATE <= NEXT_STATE;
	end if;

end if;
end process;



OUTPUT_SIGNAL_PROCESS: process(CURRENT_STATE)
begin
-- segnali default tutti a 0
LD_SHIFT_R8 <= '0';
CLEAR_R8 <= '0';
MUX_SEL_STOP_BIT <= '0';
LD_ERROR <= '0';
CLEAR_ERROR <= '0';
CLEAR_BUSY <= '0';
LD_BUSY <= '0';
LD_SHIFT_DOUT <= '0';
EN_CNT_TIME_SAMPLES <= '0';
CLEAR_CNT_TIME_SAMPLES <= '0';
EN_CNT_8_SAMPLES <= '0';
CLEAR_CNT_8_SAMPLES <= '0';
EN_CNT_SYMBOL <= '0';
CLEAR_CNT_SYMBOL <= '0';
CLEAR_DONE <= '0';
LD_DONE <= '0';
CLEAR_DOUT <= '0';
CLEAR_CNT_TIME_NOP <= '0';
EN_CNT_TIME_NOP <= '0'; 
case (CURRENT_STATE) IS
	WHEN RESET_STATE =>CLEAR_R8 <= '1';
			CLEAR_ERROR <= '1';
			CLEAR_BUSY <= '1';
			CLEAR_CNT_TIME_SAMPLES <= '1';
			CLEAR_CNT_8_SAMPLES <= '1';
			CLEAR_CNT_SYMBOL <= '1';
			CLEAR_DONE <= '1';
			CLEAR_DOUT <= '1';
			CLEAR_CNT_TIME_NOP <= '1';

	when IDLE_1 => LD_SHIFT_R8 <= '1';
			CLEAR_CNT_TIME_SAMPLES <= '1';

	when IDLE_2 => EN_CNT_TIME_SAMPLES <= '1';

	when STATE_AFTER_START_1 => LD_BUSY <= '1';
				CLEAR_DONE <= '1';
				CLEAR_ERROR <= '1';
				EN_CNT_TIME_SAMPLES <= '1';

	when STATE_AFTER_START_2 => EN_CNT_TIME_SAMPLES <= '1';

	when ANALISI_SAMPLES_START_1 => CLEAR_CNT_TIME_SAMPLES <= '1';
					EN_CNT_8_SAMPLES <= '1';
					LD_SHIFT_R8 <= '1';


	when ANALISI_SAMPLES_START_2 => EN_CNT_TIME_SAMPLES <= '1';

	when LOAD_ERROR_START => 
			CLEAR_CNT_8_SAMPLES <= '1';
			EN_CNT_TIME_NOP <= '1';
	
	when NOP_START_SYMB => EN_CNT_TIME_NOP <= '1';
	when NOP_START_SYMB_END => CLEAR_CNT_TIME_NOP <= '1';
	
	when SYMBOL_SAMPLE => LD_SHIFT_R8 <= '1';
					CLEAR_CNT_TIME_SAMPLES <= '1';
					EN_CNT_8_SAMPLES <= '1';

	when SYMBOL_WAIT => EN_CNT_TIME_SAMPLES <= '1';

	when EVALUATION_SYMBOLS => LD_SHIFT_DOUT <= '1';
					CLEAR_CNT_8_SAMPLES <= '1';
					EN_CNT_SYMBOL <= '1';

					EN_CNT_TIME_NOP <= '1';

	when NOP_SYMBOL => EN_CNT_TIME_NOP <= '1';
	when NOP_SYMBOL_END => CLEAR_CNT_TIME_NOP <= '1';



	when STOP_BIT_SAMPLES => LD_SHIFT_R8 <= '1';
					CLEAR_CNT_TIME_SAMPLES <= '1';
					EN_CNT_8_SAMPLES <= '1';

	when STOP_BIT_WAIT => EN_CNT_TIME_SAMPLES <= '1';

	when EVALUATE_ERROR_STOP => 
				CLEAR_BUSY <= '1';
				LD_DONE <= '1';
				CLEAR_CNT_TIME_SAMPLES <= '1';
				CLEAR_CNT_8_SAMPLES <= '1';
				CLEAR_CNT_SYMBOL <= '1';
				EN_CNT_TIME_SAMPLES <= '1';
				MUX_SEL_STOP_BIT <= '1';

	
	when ERROR_STOP_BIT => CLEAR_R8 <= '1';
				EN_CNT_TIME_SAMPLES <= '1';
				LD_ERROR <= '1';
	

	when MANAGE_ERROR_START_BIT => 	
					CLEAR_CNT_TIME_SAMPLES <= '1';
					CLEAR_CNT_8_SAMPLES <= '1';
					CLEAR_CNT_SYMBOL <= '1';
					CLEAR_BUSY <= '1';
					CLEAR_R8 <= '1';
					CLEAR_CNT_TIME_NOP <= '1';
					LD_ERROR <= '1';
				
				

	when OTHERS => 
			CLEAR_R8 <= '1';
			CLEAR_ERROR <= '1';
			CLEAR_BUSY <= '1';
			CLEAR_CNT_TIME_SAMPLES <= '1';
			CLEAR_CNT_8_SAMPLES <= '1';
			CLEAR_CNT_SYMBOL <= '1';
			CLEAR_DONE <= '1';
			CLEAR_DOUT <= '1';
			CLEAR_CNT_TIME_NOP <= '1';
end case;
end process;

	

	

	
	
	

	
					
	
	
			
					
			
end beh;



